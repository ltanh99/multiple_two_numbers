-- Sub Module REG:

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
 
ENTITY REG IS
PORT(
D: IN STD_LOGIC_VECTOR (7 downto 0);
CLR, ENA, CLK: IN STD_LOGIC;
Q: OUT STD_LOGIC_VECTOR (7 downto 0)
);
END REG;
 
ARCHITECTURE RTL OF REG IS
BEGIN
PROCESS(CLK, CLR)
BEGIN
IF CLR = '1' THEN
Q <= (OTHERS => '0');
ELSE
IF CLK'event and CLK = '1' THEN
IF ENA = '1' THEN
Q <= D;
ELSE null;
END IF;
END IF;
END IF;
END PROCESS;
END RTL;
