-- Module ADDER:
 
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_unsigned.all;
 
ENTITY ADDER IS
PORT(
A, B: IN STD_LOGIC_VECTOR (7 downto 0);
ENA: IN STD_LOGIC;
S: OUT STD_LOGIC_VECTOR (8 downto 0)
);
END ADDER;
 
ARCHITECTURE RTL OF ADDER IS
BEGIN
PROCESS(ENA, A, B)
BEGIN
IF ENA = '1' THEN
S <= ('0'&A)+('0'&B);
ELSE S <= '0'&A;
END IF;
END PROCESS;
END RTL;
